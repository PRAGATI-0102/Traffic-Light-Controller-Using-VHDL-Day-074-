library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TLC is

    port (
		  Clk                     : in std_logic;
		  Reset                   : in std_logic;
        State_output            : out std_logic_vector(7 downto 0));
		  
end TLC;

architecture behavioural of TLC is

	component T5 is
		
		port (
        clk : in std_logic;
        reset : in std_logic;
        T_5sec : out std_logic);
		  
	end component;
	
	component T1 is
		
		port (
        clk : in std_logic;
        reset : in std_logic;
        T_1sec : out std_logic);
		  
	end component;
	
	signal T_5sec, T_1sec : std_logic;
	--signal OUTN, OUTE, OUTS, OUTW : std_logic;

	type state is (S0,S1,S2,S3,S4,S5,S6,S7);
	
	signal Y_Present, Y_Next : state := S0;

 3	
	
	
		begin
		
		--Time Instantiation
		
		TIME1: T1 port map(clk => CLK, reset => RESET, T_1sec => T_1sec);
		TIME2: T5 port map(clk => CLK, reset => RESET, T_5sec => T_5sec);
		
		
		CLK_PROC: process (Clk,Reset)
		begin
		
			if (Clk'event and Clk = '1') then
				
				if (Reset = '1') then
				
					Y_Present <= S0;
					
				else
					
					Y_Present <= Y_Next;
				
				end if;
				
			end if;
			
			
		end process;
		
		ST_PROC: process (T_5sec, T_1sec, Y_Present)
		begin
			
			case Y_present is
				
				when S0 =>
				
					if (T_5sec = '1') then
						
						Y_Next <= S1;
						
					else
					
						Y_Next <= S0;
					
					end if;
				
				when S1 =>
				
					if (T_1sec = '1') then
						
						Y_Next <= S2;
						
					else
					
						Y_Next <= S1;
					
					end if;
						
				when S2 =>
				
					if (T_5sec = '1') then
						
						Y_Next <= S3;
						
					else
					
						Y_Next <= S2;
						
					end if;
				
				when S3 =>
				
					if (T_1sec = '1') then
						
						Y_Next <= S4;
						
					else
					
						Y_Next <= S3;
						
					end if;
				
				when S4 =>
				
					if (T_5sec = '1') then
						
						Y_Next <= S5;
						
					else
					
						Y_Next <= S4;
						
					end if;
				
				when S5 =>
				
					if (T_1sec = '1') then
						
						Y_Next <= S6;
						
					else
					
						Y_Next <= S5;
					
					end if;
				
				when S6 =>
				
					if (T_5sec = '1') then
						
						Y_Next <= S7;
						
					else
					
						Y_Next <= S6;
					
					end if;
				
				when S7 =>
				
					if (T_1sec = '1') then
						
						Y_Next <= S0;
						
					else
					
						Y_Next <= S7;
					
					end if;
						
				when others =>
				
						null;
			
			end case;
		
		end process;
		
		OUTP_PROC: process(Y_present)
		begin
		
			if (Y_present = S0) then
				State_output(7 downto 6) <= GREEN;
				State_output(5 downto 4) <= RED;
				State_output(3 downto 2) <= RED;
				State_output(1 downto 0) <= RED;
			
			elsif (Y_present = S1) then
				State_output(7 downto 6) <= YELLOW;
				State_output(5 downto 4) <= YELLOW;
				State_output(3 downto 2) <= RED;
				State_output(1 downto 0) <= RED;
				
			elsif (Y_present = S2) then
				State_output(7 downto 6) <= RED;
				State_output(5 downto 4) <= GREEN;
				State_output(3 downto 2) <= RED;
				State_output(1 downto 0) <= RED;
				
			elsif (Y_present = S3) then
				State_output(7 downto 6) <= RED;
				State_output(5 downto 4) <= YELLOW;
				State_output(3 downto 2) <= YELLOW;
				State_output(1 downto 0) <= RED;
			
			elsif (Y_present = S4) then
				State_output(7 downto 6) <= RED;
				State_output(5 downto 4) <= RED;
				State_output(3 downto 2) <= GREEN;
				State_output(1 downto 0) <= RED;
			
			elsif (Y_present = S5) then
				State_output(7 downto 6) <= RED;
				State_output(5 downto 4) <= RED;
				State_output(3 downto 2) <= YELLOW;
				State_output(1 downto 0) <= YELLOW;
			
			elsif (Y_present = S6) then
				State_output(7 downto 6) <= RED;
				State_output(5 downto 4) <= RED;
				State_output(3 downto 2) <= RED;
				State_output(1 downto 0) <= GREEN;
			
			else 
				State_output(7 downto 6) <= YELLOW;
				State_output(5 downto 4) <= RED;
				State_output(3 downto 2) <= RED;
				State_output(1 downto 0) <= YELLOW;
				
			end if;
			
		end process;

end behavioural;
